
`define FAT_COLOUR_NONEXISTENT
`define MUSCLE_COLOUR_NONEXISTENT

`define FAT_COLOUR_RAW 9'b000000000
`define MUSCLE_COLOUR_RAW 9'b000000000

`define FAT_COLOUR_RARE 9'b011000010
`define MUSCLE_COLOUR_RARE 9'b011001011

`define FAT_COLOUR_MEDIUM_RARE 9'b011111111
`define MUSCLE_COLOUR_MEDIUM_RARE 9'b100000000

`define FAT_COLOUR_MEDIUM_WELL 9'b011000111
`define MUSCLE_COLOUR_MEDIUM_WELL 9'b011111000

`define FAT_COLOUR_MEDIUM 9'b011110000
`define MUSCLE_COLOUR_MEDIUM 9'b000111000

`define FAT_COLOUR_WELL_DONE 9'b011000111
`define MUSCLE_COLOUR_WELL_DONE 9'b011110000

`define FAT_COLOUR_BURNT 9'b011111111
`define MUSCLE_COLOUR_BURNT 9'b000111111



`define x_adder0 30
`define x_adder1 70
`define x_adder2 110
`define x_adder3 30
`define x_adder4 70
`define x_adder5 110

`define y_adder0 30
`define y_adder1 30
`define y_adder2 30
`define y_adder3 70
`define y_adder4 70
`define y_adder5 70

///////////////////coordinates of fat graphics
`define x1 3
`define y1 0

`define x2 4
`define y2 0

`define x3 5
`define y3 0

`define x4 6
`define y4 0

`define x5 2
`define y5 1

`define x6 7
`define y6 1

`define x7 0
`define y7 2

`define x8 1
`define y8 2

`define x9 6
`define y9 2

`define x10 8
`define y10 2

`define x11 0
`define y11 3

`define x12 8
`define y12 3

`define x13 1
`define y13 4

`define x14 2
`define y14 4

`define x15 3
`define y15 4

`define x16 4
`define y16 4

`define x17 5
`define y17 4

`define x18 6
`define y18 4

`define x19 7
`define y19 4

`define x20 5
`define y20 5

`define x21 6
`define y21 5


/////////////////// coordinates of muscle graphics
`define q1 3
`define z1 1

`define q2 4
`define z2 1

`define q3 5
`define z3 1

`define q4 6
`define z4 1

`define q5 2
`define z5 2

`define q6 3
`define z6 2

`define q7 4
`define z7 2

`define q8 5
`define z8 2

`define q9 7
`define z9 2

`define q10 1
`define z10 3

`define q11 2
`define z11 3

`define q12 3
`define z12 3

`define q13 4
`define z13 3

`define q14 5
`define z14 3

`define q15 6
`define z15 3

`define q16 7
`define z16 3
