`define FAT_COLOUR_NONEXISTENT 9'b000000000
`define MUSCLE_COLOUR_NONEXISTENT 9'b000000000

//{66, 32, 0}
//{66, 0, 0}
`define FAT_COLOUR_RAW 9'b111000000
`define MUSCLE_COLOUR_RAW 9'b000000000

//{66, 32, 0}
//{66, 0, 0}
`define FAT_COLOUR_RARE 9'b110000000
`define MUSCLE_COLOUR_RARE 9'b000000000

//{66, 32, 0}
//{66, 0, 0}
`define FAT_COLOUR_MEDIUM_RARE 9'b101000000
`define MUSCLE_COLOUR_MEDIUM_RARE 9'b000000000

//{128, 64, 0}
//{128, 64, 64}
`define FAT_COLOUR_MEDIUM 9'b100000000
`define MUSCLE_COLOUR_MEDIUM 9'b000000000

//{128, 64, 0}
//{128, 64, 64}
`define FAT_COLOUR_MEDIUM_WELL 9'b011000000
`define MUSCLE_COLOUR_MEDIUM_WELL 9'b000000000

//{96, 32, 0}
//{96, 32, 32}
`define FAT_COLOUR_WELL_DONE 9'b010000000
`define MUSCLE_COLOUR_WELL_DONE 9'b000000000

//{66, 32, 0}
//{66, 32, 32}
// `define FAT_COLOUR_BURNT 9'b010001000
`define FAT_COLOUR_BURNT 9'b001000000
`define MUSCLE_COLOUR_BURNT 9'b000000000


//
// `define FAT_COLOUR_NONEXISTENT 9'b000000000
// `define MUSCLE_COLOUR_NONEXISTENT 9'b000000000
//
// //{66, 32, 0}
// //{66, 0, 0}
// `define FAT_COLOUR_RAW 9'b111000000
// `define MUSCLE_COLOUR_RAW 9'b000000000
//
// //{66, 32, 0}
// //{66, 0, 0}
// `define FAT_COLOUR_RARE 9'b000111000
// `define MUSCLE_COLOUR_RARE 9'b000000000
//
// //{66, 32, 0}
// //{66, 0, 0}
// `define FAT_COLOUR_MEDIUM_RARE 9'b000000111
// `define MUSCLE_COLOUR_MEDIUM_RARE 9'b000000000
//
// //{128, 64, 0}
// //{128, 64, 64}
// `define FAT_COLOUR_MEDIUM 9'b111111000
// `define MUSCLE_COLOUR_MEDIUM 9'b000000000
//
// //{128, 64, 0}
// //{128, 64, 64}
// `define FAT_COLOUR_MEDIUM_WELL 9'b111000111
// `define MUSCLE_COLOUR_MEDIUM_WELL 9'b000000000
//
// //{96, 32, 0}
// //{96, 32, 32}
// `define FAT_COLOUR_WELL_DONE 9'b000111111
// `define MUSCLE_COLOUR_WELL_DONE 9'b000000000
//
// //{66, 32, 0}
// //{66, 32, 32}
// // `define FAT_COLOUR_BURNT 9'b010001000
// `define FAT_COLOUR_BURNT 9'b111111111
// `define MUSCLE_COLOUR_BURNT 9'b000000000



`define x_adder0 30
`define x_adder1 70
`define x_adder2 110
`define x_adder3 30
`define x_adder4 70
`define x_adder5 110

`define y_adder0 30
`define y_adder1 30
`define y_adder2 30
`define y_adder3 70
`define y_adder4 70
`define y_adder5 70

///////////////////coordinates of fat graphics
`define x1 5
`define y1 0

`define x2 6
`define y2 0

`define x3 7
`define y3 0

`define x4 8
`define y4 0

`define x5 9
`define y5 0

`define x6 10
`define y6 0

`define x7 11
`define y7 0

`define x8 12
`define y8 0

`define x9 13
`define y9 0

`define x10 14
`define y10 0

`define x11 15
`define y11 0

`define x12 16
`define y12 0

`define x13 3
`define y13 1

`define x14 4
`define y14 1

`define x15 5
`define y15 1

`define x16 6
`define y16 1

`define x17 7
`define y17 1

`define x18 8
`define y18 1

`define x19 9
`define y19 1

`define x20 10
`define y20 1

`define x21 11
`define y21 1

`define x22 12
`define y22 1

`define x23 13
`define y23 1

`define x24 14
`define y24 1

`define x25 15
`define y25 1

`define x26 16
`define y26 1

`define x27 17
`define y27 1

`define x28 18
`define y28 1

`define x29 2
`define y29 2

`define x30 3
`define y30 2

`define x31 4
`define y31 2

`define x32 5
`define y32 2

`define x33 8
`define y33 2

`define x34 9
`define y34 2

`define x35 12
`define y35 2

`define x36 13
`define y36 2

`define x37 16
`define y37 2

`define x38 17
`define y38 2

`define x39 18
`define y39 2

`define x40 19
`define y40 2

`define x41 0
`define y41 3

`define x42 1
`define y42 3

`define x43 2
`define y43 3

`define x44 3
`define y44 3

`define x45 4
`define y45 3

`define x46 5
`define y46 3

`define x47 8
`define y47 3

`define x48 9
`define y48 3

`define x49 12
`define y49 3

`define x50 13
`define y50 3

`define x51 16
`define y51 3

`define x52 17
`define y52 3

`define x53 18
`define y53 3

`define x54 19
`define y54 3

`define x55 20
`define y55 3

`define x56 21
`define y56 3

`define x57 0
`define y57 4

`define x58 1
`define y58 4

`define x59 4
`define y59 4

`define x60 5
`define y60 4

`define x61 8
`define y61 4

`define x62 9
`define y62 4

`define x63 12
`define y63 4

`define x64 13
`define y64 4

`define x65 16
`define y65 4

`define x66 17
`define y66 4

`define x67 20
`define y67 4

`define x68 21
`define y68 4

`define x69 0
`define y69 5

`define x70 1
`define y70 5

`define x71 4
`define y71 5

`define x72 5
`define y72 5

`define x73 8
`define y73 5

`define x74 9
`define y74 5

`define x75 12
`define y75 5

`define x76 13
`define y76 5

`define x77 16
`define y77 5

`define x78 17
`define y78 5

`define x79 20
`define y79 5

`define x80 21
`define y80 5

`define x81 0
`define y81 6

`define x82 1
`define y82 6

`define x83 4
`define y83 6

`define x84 5
`define y84 6

`define x85 8
`define y85 6




`define x86 12
`define y86 6

`define x87 13
`define y87 6

`define x88 16
`define y88 6

`define x89 17
`define y89 6

`define x90 20
`define y90 6

`define x91 21
`define y91 6

`define x92 0
`define y92 7

`define x93 1
`define y93 7

`define x94 4
`define y94 7

`define x95 5
`define y95 7

`define x96 8
`define y96 7

`define x97 9
`define y97 7

`define x98 12
`define y98 7

`define x99 13
`define y99 7

`define x100 16
`define y100 7

`define x101 17
`define y101 7

`define x102 20
`define y102 7

`define x103 21
`define y103 7

`define x104 0
`define y104 8

`define x105 1
`define y105 8

`define x106 4
`define y106 8

`define x107 5
`define y107 8

`define x108 8
`define y108 8

`define x109 9
`define y109 8

`define x110 12
`define y110 8

`define x111 13
`define y111 8

`define x112 16
`define y112 8

`define x113 17
`define y113 8

`define x114 20
`define y114 8

`define x115 21
`define y115 8

`define x116 0
`define y116 9

`define x117 1
`define y117 9

`define x118 2
`define y118 9

`define x119 3
`define y119 9

`define x120 4
`define y120 9

`define x121 5
`define y121 9

`define x122 8
`define y122 9

`define x123 9
`define y123 9

`define x124 12
`define y124 9

`define x125 13
`define y125 9

`define x126 16
`define y126 9

`define x127 17
`define y127 9

`define x128 18
`define y128 9

`define x129 19
`define y129 9

`define x130 20
`define y130 9

`define x131 21
`define y131 9


`define x132 2
`define y132 10

`define x133 3
`define y133 10

`define x134 4
`define y134 10

`define x135 5
`define y135 10

`define x136 8
`define y136 10

`define x137 9
`define y137 10

`define x138 12
`define y138 10

`define x139 13
`define y139 10

`define x140 16
`define y140 10

`define x141 17
`define y141 10

`define x142 18
`define y142 10

`define x143 19
`define y143 10


`define x144 3
`define y144 11

`define x145 4
`define y145 11

`define x146 5
`define y146 11

`define x147 6
`define y147 11

`define x148 7
`define y148 11

`define x149 8
`define y149 11

`define x150 9
`define y150 11

`define x151 10
`define y151 11

`define x152 11
`define y152 11

`define x153 12
`define y153 11

`define x154 13
`define y154 11

`define x155 14
`define y155 11

`define x156 15
`define y156 11

`define x157 16
`define y157 11

`define x158 17
`define y158 11

`define x159 18
`define y159 11

`define x160 5
`define y160 12

`define x161 6
`define y161 12

`define x162 7
`define y162 12

`define x163 8
`define y163 12

`define x164 9
`define y164 12

`define x165 10
`define y165 12

`define x166 11
`define y166 12

`define x167 12
`define y167 12

`define x168 13
`define y168 12

`define x169 14
`define y169 12

`define x170 15
`define y170 12

`define x171 16
`define y171 12

`define x172 9
`define y172 6


/////////////////// coordinates of muscle graphics
`define q1 6
`define z1 2

`define q2 7
`define z2 2

`define q3 10
`define z3 2

`define q4 11
`define z4 2

`define q5 14
`define z5 2

`define q6 15
`define z6 2

`define q7 6
`define z7 3

`define q8 7
`define z8 3

`define q9 10
`define z9 3

`define q10 11
`define z10 3

`define q11 14
`define z11 3

`define q12 15
`define z12 3

`define q13 2
`define z13 4

`define q14 3
`define z14 4

`define q15 6
`define z15 4

`define q16 7
`define z16 4

`define q17 10
`define z17 4

`define q18 11
`define z18 4

`define q19 14
`define z19 4

`define q20 15
`define z20 4

`define q21 18
`define z21 4

`define q22 19
`define z22 4

`define q23 2
`define z23 5

`define q24 3
`define z24 5

`define q25 6
`define z25 5

`define q26 7
`define z26 5

`define q27 10
`define z27 5

`define q28 11
`define z28 5

`define q29 14
`define z29 5

`define q30 15
`define z30 5

`define q31 18
`define z31 5

`define q32 19
`define z32 5

`define q33 2
`define z33 6

`define q34 3
`define z34 6

`define q35 6
`define z35 6

`define q36 7
`define z36 6

`define q37 10
`define z37 6

`define q38 11
`define z38 6

`define q39 14
`define z39 6

`define q40 15
`define z40 6

`define q41 18
`define z41 6

`define q42 19
`define z42 6

`define q43 2
`define z43 7

`define q44 3
`define z44 7

`define q45 6
`define z45 7

`define q46 7
`define z46 7

`define q47 10
`define z47 7

`define q48 11
`define z48 7

`define q49 14
`define z49 7

`define q50 15
`define z50 7

`define q51 18
`define z51 7

`define q52 19
`define z52 7

`define q53 2
`define z53 8

`define q54 3
`define z54 8

`define q55 6
`define z55 8

`define q56 7
`define z56 8

`define q57 10
`define z57 8

`define q58 11
`define z58 8

`define q59 14
`define z59 8

`define q60 15
`define z60 8

`define q61 18
`define z61 8

`define q62 19
`define z62 8


`define q63 6
`define z63 9

`define q64 7
`define z64 9

`define q65 10
`define z65 9

`define q66 11
`define z66 9

`define q67 14
`define z67 9

`define q68 15
`define z68 9


`define q69 6
`define z69 10

`define q70 7
`define z70 10

`define q71 10
`define z71 10

`define q72 11
`define z72 10

`define q73 14
`define z73 10

`define q74 15
`define z74 10
